module fdiv(
    input  logic clk,rst,
    input  logic [31:0] x,y,
    output logic [31:0] z
);
    logic [35:0] init_grad [1023:0];
    logic xs,ys;
    logic [7:0] xe,ye;
    logic [23:0] xm;
    logic [9:0]  key;
    logic [12:0] diff;
    assign {xs, xe, xm[22:0]} = x;
    assign xm[23] = 1'b1;
    assign {ys, ye, key, diff} = y;
    logic unsigned [34:0] init;
    logic unsigned [12:0] grad;
    assign init = {init_grad[key][35:13], 12'b0} ;
    assign grad = init_grad[key][12:0];
    logic unsigned [35:0] ym_;
    assign ym_ = init - diff * grad;
    logic [23:0] ym;
    assign ym  = {1'b1, ym_[34:12]};
    logic [47:0] m_;
    assign m_ = xm * ym;
    logic [22:0] m;
    assign m = m_[47] ? m_[46:24] : m_[45:23];
    logic s;
    assign s = xs ^ ys;

    logic [8:0] e_;
    assign e_  = {1'b0, xe} - {1'b0, ye} + 9'd126;
    logic [8:0] e_p1 ;
    assign e_p1 = e_ + 1;

    logic [7:0] e;
    assign e = m_[47] ? e_p1[7:0] : e_[7:0];
    assign z = {s,e,m};



    initial begin
        
init_grad[ 0 ] = 36'hfffffbff7 ;
init_grad[ 1 ] = 36'hff801bfe8 ;
init_grad[ 2 ] = 36'hff007bfd8 ;
init_grad[ 3 ] = 36'hfe8119fc8 ;
init_grad[ 4 ] = 36'hfe01f9fb8 ;
init_grad[ 5 ] = 36'hfd8317fa8 ;
init_grad[ 6 ] = 36'hfd0475f98 ;
init_grad[ 7 ] = 36'hfc8611f89 ;
init_grad[ 8 ] = 36'hfc07ebf79 ;
init_grad[ 9 ] = 36'hfb8a05f6a ;
init_grad[ 10 ] = 36'hfb0c5bf5a ;
init_grad[ 11 ] = 36'hfa8ef1f4b ;
init_grad[ 12 ] = 36'hfa11c5f3b ;
init_grad[ 13 ] = 36'hf994d7f2c ;
init_grad[ 14 ] = 36'hf91827f1c ;
init_grad[ 15 ] = 36'hf89bb3f0d ;
init_grad[ 16 ] = 36'hf81f7defe ;
init_grad[ 17 ] = 36'hf7a383eef ;
init_grad[ 18 ] = 36'hf727c7edf ;
init_grad[ 19 ] = 36'hf6ac49ed0 ;
init_grad[ 20 ] = 36'hf63105ec1 ;
init_grad[ 21 ] = 36'hf5b5ffeb2 ;
init_grad[ 22 ] = 36'hf53b35ea3 ;
init_grad[ 23 ] = 36'hf4c0a7e94 ;
init_grad[ 24 ] = 36'hf44655e85 ;
init_grad[ 25 ] = 36'hf3cc3fe76 ;
init_grad[ 26 ] = 36'hf35263e67 ;
init_grad[ 27 ] = 36'hf2d8c3e59 ;
init_grad[ 28 ] = 36'hf25f5fe4a ;
init_grad[ 29 ] = 36'hf1e635e3b ;
init_grad[ 30 ] = 36'hf16d47e2c ;
init_grad[ 31 ] = 36'hf0f493e1e ;
init_grad[ 32 ] = 36'hf07c1be0f ;
init_grad[ 33 ] = 36'hf003dbe01 ;
init_grad[ 34 ] = 36'hef8bd7df2 ;
init_grad[ 35 ] = 36'hef140bde4 ;
init_grad[ 36 ] = 36'hee9c7bdd5 ;
init_grad[ 37 ] = 36'hee2523dc7 ;
init_grad[ 38 ] = 36'hedae05db9 ;
init_grad[ 39 ] = 36'hed3721daa ;
init_grad[ 40 ] = 36'hecc077d9c ;
init_grad[ 41 ] = 36'hec4a05d8e ;
init_grad[ 42 ] = 36'hebd3cbd80 ;
init_grad[ 43 ] = 36'heb5dcbd71 ;
init_grad[ 44 ] = 36'heae803d63 ;
init_grad[ 45 ] = 36'hea7273d55 ;
init_grad[ 46 ] = 36'he9fd1dd47 ;
init_grad[ 47 ] = 36'he987fdd39 ;
init_grad[ 48 ] = 36'he91317d2b ;
init_grad[ 49 ] = 36'he89e67d1d ;
init_grad[ 50 ] = 36'he829efd10 ;
init_grad[ 51 ] = 36'he7b5afd02 ;
init_grad[ 52 ] = 36'he741a5cf4 ;
init_grad[ 53 ] = 36'he6cdd3ce6 ;
init_grad[ 54 ] = 36'he65a39cd8 ;
init_grad[ 55 ] = 36'he5e6d5ccb ;
init_grad[ 56 ] = 36'he573a9cbd ;
init_grad[ 57 ] = 36'he500b1cb0 ;
init_grad[ 58 ] = 36'he48df1ca2 ;
init_grad[ 59 ] = 36'he41b67c94 ;
init_grad[ 60 ] = 36'he3a913c87 ;
init_grad[ 61 ] = 36'he336f5c7a ;
init_grad[ 62 ] = 36'he2c50dc6c ;
init_grad[ 63 ] = 36'he2535bc5f ;
init_grad[ 64 ] = 36'he1e1ddc51 ;
init_grad[ 65 ] = 36'he17095c44 ;
init_grad[ 66 ] = 36'he0ff83c37 ;
init_grad[ 67 ] = 36'he08ea5c2a ;
init_grad[ 68 ] = 36'he01dfdc1c ;
init_grad[ 69 ] = 36'hdfad89c0f ;
init_grad[ 70 ] = 36'hdf3d4bc02 ;
init_grad[ 71 ] = 36'hdecd41bf5 ;
init_grad[ 72 ] = 36'hde5d69be8 ;
init_grad[ 73 ] = 36'hddedc7bdb ;
init_grad[ 74 ] = 36'hdd7e59bce ;
init_grad[ 75 ] = 36'hdd0f1fbc1 ;
init_grad[ 76 ] = 36'hdca019bb4 ;
init_grad[ 77 ] = 36'hdc3147ba7 ;
init_grad[ 78 ] = 36'hdbc2a7b9a ;
init_grad[ 79 ] = 36'hdb543bb8e ;
init_grad[ 80 ] = 36'hdae603b81 ;
init_grad[ 81 ] = 36'hda77fdb74 ;
init_grad[ 82 ] = 36'hda0a2bb67 ;
init_grad[ 83 ] = 36'hd99c8bb5b ;
init_grad[ 84 ] = 36'hd92f1db4e ;
init_grad[ 85 ] = 36'hd8c1e3b42 ;
init_grad[ 86 ] = 36'hd854dbb35 ;
init_grad[ 87 ] = 36'hd7e805b28 ;
init_grad[ 88 ] = 36'hd77b61b1c ;
init_grad[ 89 ] = 36'hd70eefb10 ;
init_grad[ 90 ] = 36'hd6a2afb03 ;
init_grad[ 91 ] = 36'hd636a1af7 ;
init_grad[ 92 ] = 36'hd5cac3aea ;
init_grad[ 93 ] = 36'hd55f19ade ;
init_grad[ 94 ] = 36'hd4f39fad2 ;
init_grad[ 95 ] = 36'hd48855ac5 ;
init_grad[ 96 ] = 36'hd41d3dab9 ;
init_grad[ 97 ] = 36'hd3b257aad ;
init_grad[ 98 ] = 36'hd347a1aa1 ;
init_grad[ 99 ] = 36'hd2dd1ba95 ;
init_grad[ 100 ] = 36'hd272c7a89 ;
init_grad[ 101 ] = 36'hd208a1a7d ;
init_grad[ 102 ] = 36'hd19eada71 ;
init_grad[ 103 ] = 36'hd134e9a65 ;
init_grad[ 104 ] = 36'hd0cb55a59 ;
init_grad[ 105 ] = 36'hd061f1a4d ;
init_grad[ 106 ] = 36'hcff8bda41 ;
init_grad[ 107 ] = 36'hcf8fb7a35 ;
init_grad[ 108 ] = 36'hcf26e1a29 ;
init_grad[ 109 ] = 36'hcebe3ba1d ;
init_grad[ 110 ] = 36'hce55c5a11 ;
init_grad[ 111 ] = 36'hcded7da06 ;
init_grad[ 112 ] = 36'hcd85659fa ;
init_grad[ 113 ] = 36'hcd1d7b9ee ;
init_grad[ 114 ] = 36'hccb5bf9e3 ;
init_grad[ 115 ] = 36'hcc4e339d7 ;
init_grad[ 116 ] = 36'hcbe6d59cb ;
init_grad[ 117 ] = 36'hcb7fa59c0 ;
init_grad[ 118 ] = 36'hcb18a59b4 ;
init_grad[ 119 ] = 36'hcab1d19a9 ;
init_grad[ 120 ] = 36'hca4b2d99d ;
init_grad[ 121 ] = 36'hc9e4b5992 ;
init_grad[ 122 ] = 36'hc97e6b986 ;
init_grad[ 123 ] = 36'hc9185197b ;
init_grad[ 124 ] = 36'hc8b261970 ;
init_grad[ 125 ] = 36'hc84ca1964 ;
init_grad[ 126 ] = 36'hc7e70d959 ;
init_grad[ 127 ] = 36'hc781a794e ;
init_grad[ 128 ] = 36'hc71c6f943 ;
init_grad[ 129 ] = 36'hc6b761937 ;
init_grad[ 130 ] = 36'hc6528392c ;
init_grad[ 131 ] = 36'hc5edcf921 ;
init_grad[ 132 ] = 36'hc58949916 ;
init_grad[ 133 ] = 36'hc524ef90b ;
init_grad[ 134 ] = 36'hc4c0c3900 ;
init_grad[ 135 ] = 36'hc45cc18f5 ;
init_grad[ 136 ] = 36'hc3f8ed8ea ;
init_grad[ 137 ] = 36'hc395438df ;
init_grad[ 138 ] = 36'hc331c78d4 ;
init_grad[ 139 ] = 36'hc2ce758c9 ;
init_grad[ 140 ] = 36'hc26b4f8be ;
init_grad[ 141 ] = 36'hc208578b3 ;
init_grad[ 142 ] = 36'hc1a5878a8 ;
init_grad[ 143 ] = 36'hc142e589d ;
init_grad[ 144 ] = 36'hc0e06d893 ;
init_grad[ 145 ] = 36'hc07e1f888 ;
init_grad[ 146 ] = 36'hc01bff87d ;
init_grad[ 147 ] = 36'hbfba07873 ;
init_grad[ 148 ] = 36'hbf583b868 ;
init_grad[ 149 ] = 36'hbef69b85d ;
init_grad[ 150 ] = 36'hbe9523853 ;
init_grad[ 151 ] = 36'hbe33d7848 ;
init_grad[ 152 ] = 36'hbdd2b583d ;
init_grad[ 153 ] = 36'hbd71bd833 ;
init_grad[ 154 ] = 36'hbd10ef828 ;
init_grad[ 155 ] = 36'hbcb04d81e ;
init_grad[ 156 ] = 36'hbc4fd3813 ;
init_grad[ 157 ] = 36'hbbef83809 ;
init_grad[ 158 ] = 36'hbb8f5d7ff ;
init_grad[ 159 ] = 36'hbb2f617f4 ;
init_grad[ 160 ] = 36'hbacf8d7ea ;
init_grad[ 161 ] = 36'hba6fe57e0 ;
init_grad[ 162 ] = 36'hba10657d5 ;
init_grad[ 163 ] = 36'hb9b10d7cb ;
init_grad[ 164 ] = 36'hb951df7c1 ;
init_grad[ 165 ] = 36'hb8f2db7b7 ;
init_grad[ 166 ] = 36'hb893ff7ac ;
init_grad[ 167 ] = 36'hb8354b7a2 ;
init_grad[ 168 ] = 36'hb7d6c1798 ;
init_grad[ 169 ] = 36'hb7785f78e ;
init_grad[ 170 ] = 36'hb71a25784 ;
init_grad[ 171 ] = 36'hb6bc1377a ;
init_grad[ 172 ] = 36'hb65e2b770 ;
init_grad[ 173 ] = 36'hb6006b766 ;
init_grad[ 174 ] = 36'hb5a2d175c ;
init_grad[ 175 ] = 36'hb54561752 ;
init_grad[ 176 ] = 36'hb4e817748 ;
init_grad[ 177 ] = 36'hb48af773e ;
init_grad[ 178 ] = 36'hb42dfd734 ;
init_grad[ 179 ] = 36'hb3d12b72a ;
init_grad[ 180 ] = 36'hb37481720 ;
init_grad[ 181 ] = 36'hb317ff716 ;
init_grad[ 182 ] = 36'hb2bba370d ;
init_grad[ 183 ] = 36'hb25f6f703 ;
init_grad[ 184 ] = 36'hb203616f9 ;
init_grad[ 185 ] = 36'hb1a77b6ef ;
init_grad[ 186 ] = 36'hb14bbb6e6 ;
init_grad[ 187 ] = 36'hb0f0216dc ;
init_grad[ 188 ] = 36'hb094af6d2 ;
init_grad[ 189 ] = 36'hb039656c9 ;
init_grad[ 190 ] = 36'hafde3f6bf ;
init_grad[ 191 ] = 36'haf83416b6 ;
init_grad[ 192 ] = 36'haf28696ac ;
init_grad[ 193 ] = 36'haecdb76a2 ;
init_grad[ 194 ] = 36'hae732b699 ;
init_grad[ 195 ] = 36'hae18c568f ;
init_grad[ 196 ] = 36'hadbe85686 ;
init_grad[ 197 ] = 36'had646b67d ;
init_grad[ 198 ] = 36'had0a77673 ;
init_grad[ 199 ] = 36'hacb0a766a ;
init_grad[ 200 ] = 36'hac56ff660 ;
init_grad[ 201 ] = 36'habfd7b657 ;
init_grad[ 202 ] = 36'haba41d64e ;
init_grad[ 203 ] = 36'hab4ae3644 ;
init_grad[ 204 ] = 36'haaf1cf63b ;
init_grad[ 205 ] = 36'haa98e1632 ;
init_grad[ 206 ] = 36'haa4017629 ;
init_grad[ 207 ] = 36'ha9e77361f ;
init_grad[ 208 ] = 36'ha98ef3616 ;
init_grad[ 209 ] = 36'ha9369760d ;
init_grad[ 210 ] = 36'ha8de61604 ;
init_grad[ 211 ] = 36'ha8864f5fb ;
init_grad[ 212 ] = 36'ha82e635f2 ;
init_grad[ 213 ] = 36'ha7d6995e9 ;
init_grad[ 214 ] = 36'ha77ef55e0 ;
init_grad[ 215 ] = 36'ha727735d7 ;
init_grad[ 216 ] = 36'ha6d0175ce ;
init_grad[ 217 ] = 36'ha678df5c5 ;
init_grad[ 218 ] = 36'ha621cb5bc ;
init_grad[ 219 ] = 36'ha5cadb5b3 ;
init_grad[ 220 ] = 36'ha5740d5aa ;
init_grad[ 221 ] = 36'ha51d655a1 ;
init_grad[ 222 ] = 36'ha4c6df598 ;
init_grad[ 223 ] = 36'ha4707d58f ;
init_grad[ 224 ] = 36'ha41a3f586 ;
init_grad[ 225 ] = 36'ha3c42357d ;
init_grad[ 226 ] = 36'ha36e2b575 ;
init_grad[ 227 ] = 36'ha3185756c ;
init_grad[ 228 ] = 36'ha2c2a5563 ;
init_grad[ 229 ] = 36'ha26d1755a ;
init_grad[ 230 ] = 36'ha217ab552 ;
init_grad[ 231 ] = 36'ha1c263549 ;
init_grad[ 232 ] = 36'ha16d3d540 ;
init_grad[ 233 ] = 36'ha11839538 ;
init_grad[ 234 ] = 36'ha0c35952f ;
init_grad[ 235 ] = 36'ha06e9b526 ;
init_grad[ 236 ] = 36'ha019ff51e ;
init_grad[ 237 ] = 36'h9fc585515 ;
init_grad[ 238 ] = 36'h9f712f50d ;
init_grad[ 239 ] = 36'h9f1cf9504 ;
init_grad[ 240 ] = 36'h9ec8e74fc ;
init_grad[ 241 ] = 36'h9e74f54f3 ;
init_grad[ 242 ] = 36'h9e21274eb ;
init_grad[ 243 ] = 36'h9dcd794e2 ;
init_grad[ 244 ] = 36'h9d79ef4da ;
init_grad[ 245 ] = 36'h9d26854d1 ;
init_grad[ 246 ] = 36'h9cd33d4c9 ;
init_grad[ 247 ] = 36'h9c80174c1 ;
init_grad[ 248 ] = 36'h9c2d134b8 ;
init_grad[ 249 ] = 36'h9bda2f4b0 ;
init_grad[ 250 ] = 36'h9b876d4a8 ;
init_grad[ 251 ] = 36'h9b34cb49f ;
init_grad[ 252 ] = 36'h9ae24b497 ;
init_grad[ 253 ] = 36'h9a8fed48f ;
init_grad[ 254 ] = 36'h9a3daf487 ;
init_grad[ 255 ] = 36'h99eb9347e ;
init_grad[ 256 ] = 36'h999997476 ;
init_grad[ 257 ] = 36'h9947bb46e ;
init_grad[ 258 ] = 36'h98f601466 ;
init_grad[ 259 ] = 36'h98a46745e ;
init_grad[ 260 ] = 36'h9852ef456 ;
init_grad[ 261 ] = 36'h98019544e ;
init_grad[ 262 ] = 36'h97b05d446 ;
init_grad[ 263 ] = 36'h975f4543d ;
init_grad[ 264 ] = 36'h970e4d435 ;
init_grad[ 265 ] = 36'h96bd7542d ;
init_grad[ 266 ] = 36'h966cbd425 ;
init_grad[ 267 ] = 36'h961c2541d ;
init_grad[ 268 ] = 36'h95cbaf415 ;
init_grad[ 269 ] = 36'h957b5740e ;
init_grad[ 270 ] = 36'h952b1f406 ;
init_grad[ 271 ] = 36'h94db053fe ;
init_grad[ 272 ] = 36'h948b0d3f6 ;
init_grad[ 273 ] = 36'h943b353ee ;
init_grad[ 274 ] = 36'h93eb7b3e6 ;
init_grad[ 275 ] = 36'h939be13de ;
init_grad[ 276 ] = 36'h934c653d6 ;
init_grad[ 277 ] = 36'h92fd093cf ;
init_grad[ 278 ] = 36'h92adcd3c7 ;
init_grad[ 279 ] = 36'h925eb13bf ;
init_grad[ 280 ] = 36'h920fb33b7 ;
init_grad[ 281 ] = 36'h91c0d33b0 ;
init_grad[ 282 ] = 36'h9172133a8 ;
init_grad[ 283 ] = 36'h9123713a0 ;
init_grad[ 284 ] = 36'h90d4ef398 ;
init_grad[ 285 ] = 36'h90868b391 ;
init_grad[ 286 ] = 36'h903845389 ;
init_grad[ 287 ] = 36'h8fea1f382 ;
init_grad[ 288 ] = 36'h8f9c1737a ;
init_grad[ 289 ] = 36'h8f4e2d372 ;
init_grad[ 290 ] = 36'h8f006136b ;
init_grad[ 291 ] = 36'h8eb2b5363 ;
init_grad[ 292 ] = 36'h8e652535c ;
init_grad[ 293 ] = 36'h8e17b5354 ;
init_grad[ 294 ] = 36'h8dca6134d ;
init_grad[ 295 ] = 36'h8d7d2d345 ;
init_grad[ 296 ] = 36'h8d301733e ;
init_grad[ 297 ] = 36'h8ce31d336 ;
init_grad[ 298 ] = 36'h8c964332f ;
init_grad[ 299 ] = 36'h8c4985327 ;
init_grad[ 300 ] = 36'h8bfce5320 ;
init_grad[ 301 ] = 36'h8bb063319 ;
init_grad[ 302 ] = 36'h8b63ff311 ;
init_grad[ 303 ] = 36'h8b17b930a ;
init_grad[ 304 ] = 36'h8acb8f303 ;
init_grad[ 305 ] = 36'h8a7f832fb ;
init_grad[ 306 ] = 36'h8a33932f4 ;
init_grad[ 307 ] = 36'h89e7c12ed ;
init_grad[ 308 ] = 36'h899c0d2e5 ;
init_grad[ 309 ] = 36'h8950752de ;
init_grad[ 310 ] = 36'h8904fb2d7 ;
init_grad[ 311 ] = 36'h88b99d2d0 ;
init_grad[ 312 ] = 36'h886e5d2c8 ;
init_grad[ 313 ] = 36'h8823392c1 ;
init_grad[ 314 ] = 36'h87d8312ba ;
init_grad[ 315 ] = 36'h878d472b3 ;
init_grad[ 316 ] = 36'h8742792ac ;
init_grad[ 317 ] = 36'h86f7c92a5 ;
init_grad[ 318 ] = 36'h86ad3329e ;
init_grad[ 319 ] = 36'h8662bb296 ;
init_grad[ 320 ] = 36'h86185f28f ;
init_grad[ 321 ] = 36'h85ce1f288 ;
init_grad[ 322 ] = 36'h8583fd281 ;
init_grad[ 323 ] = 36'h8539f527a ;
init_grad[ 324 ] = 36'h84f009273 ;
init_grad[ 325 ] = 36'h84a63b26c ;
init_grad[ 326 ] = 36'h845c87265 ;
init_grad[ 327 ] = 36'h8412f125e ;
init_grad[ 328 ] = 36'h83c975257 ;
init_grad[ 329 ] = 36'h838015250 ;
init_grad[ 330 ] = 36'h8336d324a ;
init_grad[ 331 ] = 36'h82edab243 ;
init_grad[ 332 ] = 36'h82a49d23c ;
init_grad[ 333 ] = 36'h825bad235 ;
init_grad[ 334 ] = 36'h8212d722e ;
init_grad[ 335 ] = 36'h81ca1d227 ;
init_grad[ 336 ] = 36'h81817f220 ;
init_grad[ 337 ] = 36'h8138fd219 ;
init_grad[ 338 ] = 36'h80f095213 ;
init_grad[ 339 ] = 36'h80a84720c ;
init_grad[ 340 ] = 36'h806015205 ;
init_grad[ 341 ] = 36'h8017ff1fe ;
init_grad[ 342 ] = 36'h7fd0031f8 ;
init_grad[ 343 ] = 36'h7f88231f1 ;
init_grad[ 344 ] = 36'h7f405d1ea ;
init_grad[ 345 ] = 36'h7ef8b31e4 ;
init_grad[ 346 ] = 36'h7eb1231dd ;
init_grad[ 347 ] = 36'h7e69ad1d6 ;
init_grad[ 348 ] = 36'h7e22531d0 ;
init_grad[ 349 ] = 36'h7ddb131c9 ;
init_grad[ 350 ] = 36'h7d93ed1c2 ;
init_grad[ 351 ] = 36'h7d4ce31bc ;
init_grad[ 352 ] = 36'h7d05f11b5 ;
init_grad[ 353 ] = 36'h7cbf1b1ae ;
init_grad[ 354 ] = 36'h7c785f1a8 ;
init_grad[ 355 ] = 36'h7c31bf1a1 ;
init_grad[ 356 ] = 36'h7beb3719b ;
init_grad[ 357 ] = 36'h7ba4c9194 ;
init_grad[ 358 ] = 36'h7b5e7718e ;
init_grad[ 359 ] = 36'h7b183d187 ;
init_grad[ 360 ] = 36'h7ad21f181 ;
init_grad[ 361 ] = 36'h7a8c1917a ;
init_grad[ 362 ] = 36'h7a462d174 ;
init_grad[ 363 ] = 36'h7a005d16d ;
init_grad[ 364 ] = 36'h79baa5167 ;
init_grad[ 365 ] = 36'h797507161 ;
init_grad[ 366 ] = 36'h792f8315a ;
init_grad[ 367 ] = 36'h78ea17154 ;
init_grad[ 368 ] = 36'h78a4c514d ;
init_grad[ 369 ] = 36'h785f8f147 ;
init_grad[ 370 ] = 36'h781a6f141 ;
init_grad[ 371 ] = 36'h77d56b13a ;
init_grad[ 372 ] = 36'h77907f134 ;
init_grad[ 373 ] = 36'h774bad12e ;
init_grad[ 374 ] = 36'h7706f3128 ;
init_grad[ 375 ] = 36'h76c253121 ;
init_grad[ 376 ] = 36'h767dcd11b ;
init_grad[ 377 ] = 36'h76395f115 ;
init_grad[ 378 ] = 36'h75f50910f ;
init_grad[ 379 ] = 36'h75b0cd108 ;
init_grad[ 380 ] = 36'h756cab102 ;
init_grad[ 381 ] = 36'h75289f0fc ;
init_grad[ 382 ] = 36'h74e4af0f6 ;
init_grad[ 383 ] = 36'h74a0d50f0 ;
init_grad[ 384 ] = 36'h745d150e9 ;
init_grad[ 385 ] = 36'h74196d0e3 ;
init_grad[ 386 ] = 36'h73d5df0dd ;
init_grad[ 387 ] = 36'h7392690d7 ;
init_grad[ 388 ] = 36'h734f0b0d1 ;
init_grad[ 389 ] = 36'h730bc50cb ;
init_grad[ 390 ] = 36'h72c8970c5 ;
init_grad[ 391 ] = 36'h7285830bf ;
init_grad[ 392 ] = 36'h7242850b9 ;
init_grad[ 393 ] = 36'h71ffa10b3 ;
init_grad[ 394 ] = 36'h71bcd50ad ;
init_grad[ 395 ] = 36'h717a210a7 ;
init_grad[ 396 ] = 36'h7137850a1 ;
init_grad[ 397 ] = 36'h70f50109b ;
init_grad[ 398 ] = 36'h70b295095 ;
init_grad[ 399 ] = 36'h70704108f ;
init_grad[ 400 ] = 36'h702e03089 ;
init_grad[ 401 ] = 36'h6febdf083 ;
init_grad[ 402 ] = 36'h6fa9d307d ;
init_grad[ 403 ] = 36'h6f67dd077 ;
init_grad[ 404 ] = 36'h6f25ff071 ;
init_grad[ 405 ] = 36'h6ee43906b ;
init_grad[ 406 ] = 36'h6ea28b065 ;
init_grad[ 407 ] = 36'h6e60f505f ;
init_grad[ 408 ] = 36'h6e1f7505a ;
init_grad[ 409 ] = 36'h6dde0d054 ;
init_grad[ 410 ] = 36'h6d9cbd04e ;
init_grad[ 411 ] = 36'h6d5b83048 ;
init_grad[ 412 ] = 36'h6d1a61042 ;
init_grad[ 413 ] = 36'h6cd95503c ;
init_grad[ 414 ] = 36'h6c9861037 ;
init_grad[ 415 ] = 36'h6c5785031 ;
init_grad[ 416 ] = 36'h6c16bf02b ;
init_grad[ 417 ] = 36'h6bd611025 ;
init_grad[ 418 ] = 36'h6b9579020 ;
init_grad[ 419 ] = 36'h6b54f901a ;
init_grad[ 420 ] = 36'h6b148f014 ;
init_grad[ 421 ] = 36'h6ad43b00f ;
init_grad[ 422 ] = 36'h6a93ff009 ;
init_grad[ 423 ] = 36'h6a53d9003 ;
init_grad[ 424 ] = 36'h6a13caffd ;
init_grad[ 425 ] = 36'h69d3d2ff8 ;
init_grad[ 426 ] = 36'h6993f0ff2 ;
init_grad[ 427 ] = 36'h695426fed ;
init_grad[ 428 ] = 36'h691470fe7 ;
init_grad[ 429 ] = 36'h68d4d2fe1 ;
init_grad[ 430 ] = 36'h68954afdc ;
init_grad[ 431 ] = 36'h6855dafd6 ;
init_grad[ 432 ] = 36'h68167efd1 ;
init_grad[ 433 ] = 36'h67d73afcb ;
init_grad[ 434 ] = 36'h67980cfc6 ;
init_grad[ 435 ] = 36'h6758f2fc0 ;
init_grad[ 436 ] = 36'h6719f0fbb ;
init_grad[ 437 ] = 36'h66db04fb5 ;
init_grad[ 438 ] = 36'h669c2efb0 ;
init_grad[ 439 ] = 36'h665d6efaa ;
init_grad[ 440 ] = 36'h661ec4fa5 ;
init_grad[ 441 ] = 36'h65e030f9f ;
init_grad[ 442 ] = 36'h65a1b2f9a ;
init_grad[ 443 ] = 36'h656348f94 ;
init_grad[ 444 ] = 36'h6524f6f8f ;
init_grad[ 445 ] = 36'h64e6b8f89 ;
init_grad[ 446 ] = 36'h64a890f84 ;
init_grad[ 447 ] = 36'h646a80f7f ;
init_grad[ 448 ] = 36'h642c82f79 ;
init_grad[ 449 ] = 36'h63ee9cf74 ;
init_grad[ 450 ] = 36'h63b0caf6e ;
init_grad[ 451 ] = 36'h637310f69 ;
init_grad[ 452 ] = 36'h633568f64 ;
init_grad[ 453 ] = 36'h62f7d8f5e ;
init_grad[ 454 ] = 36'h62ba5cf59 ;
init_grad[ 455 ] = 36'h627cf6f54 ;
init_grad[ 456 ] = 36'h623fa4f4e ;
init_grad[ 457 ] = 36'h620268f49 ;
init_grad[ 458 ] = 36'h61c542f44 ;
init_grad[ 459 ] = 36'h618830f3f ;
init_grad[ 460 ] = 36'h614b34f39 ;
init_grad[ 461 ] = 36'h610e4cf34 ;
init_grad[ 462 ] = 36'h60d17af2f ;
init_grad[ 463 ] = 36'h6094bcf2a ;
init_grad[ 464 ] = 36'h605814f24 ;
init_grad[ 465 ] = 36'h601b80f1f ;
init_grad[ 466 ] = 36'h5fdf00f1a ;
init_grad[ 467 ] = 36'h5fa296f15 ;
init_grad[ 468 ] = 36'h5f6640f10 ;
init_grad[ 469 ] = 36'h5f2a00f0b ;
init_grad[ 470 ] = 36'h5eedd4f05 ;
init_grad[ 471 ] = 36'h5eb1bcf00 ;
init_grad[ 472 ] = 36'h5e75b8efb ;
init_grad[ 473 ] = 36'h5e39caef6 ;
init_grad[ 474 ] = 36'h5dfdf0ef1 ;
init_grad[ 475 ] = 36'h5dc22aeec ;
init_grad[ 476 ] = 36'h5d867aee7 ;
init_grad[ 477 ] = 36'h5d4adcee2 ;
init_grad[ 478 ] = 36'h5d0f54edd ;
init_grad[ 479 ] = 36'h5cd3e0ed7 ;
init_grad[ 480 ] = 36'h5c9880ed2 ;
init_grad[ 481 ] = 36'h5c5d34ecd ;
init_grad[ 482 ] = 36'h5c21fcec8 ;
init_grad[ 483 ] = 36'h5be6daec3 ;
init_grad[ 484 ] = 36'h5babcaebe ;
init_grad[ 485 ] = 36'h5b70ceeb9 ;
init_grad[ 486 ] = 36'h5b35e6eb4 ;
init_grad[ 487 ] = 36'h5afb14eaf ;
init_grad[ 488 ] = 36'h5ac054eaa ;
init_grad[ 489 ] = 36'h5a85a8ea5 ;
init_grad[ 490 ] = 36'h5a4b10ea0 ;
init_grad[ 491 ] = 36'h5a108ce9c ;
init_grad[ 492 ] = 36'h59d61ce97 ;
init_grad[ 493 ] = 36'h599bc0e92 ;
init_grad[ 494 ] = 36'h596178e8d ;
init_grad[ 495 ] = 36'h592742e88 ;
init_grad[ 496 ] = 36'h58ed20e83 ;
init_grad[ 497 ] = 36'h58b312e7e ;
init_grad[ 498 ] = 36'h587918e79 ;
init_grad[ 499 ] = 36'h583f30e74 ;
init_grad[ 500 ] = 36'h58055ee70 ;
init_grad[ 501 ] = 36'h57cb9ee6b ;
init_grad[ 502 ] = 36'h5791f0e66 ;
init_grad[ 503 ] = 36'h575858e61 ;
init_grad[ 504 ] = 36'h571ed2e5c ;
init_grad[ 505 ] = 36'h56e55ee57 ;
init_grad[ 506 ] = 36'h56abfee53 ;
init_grad[ 507 ] = 36'h5672b2e4e ;
init_grad[ 508 ] = 36'h56397ae49 ;
init_grad[ 509 ] = 36'h560052e44 ;
init_grad[ 510 ] = 36'h55c740e40 ;
init_grad[ 511 ] = 36'h558e40e3b ;
init_grad[ 512 ] = 36'h555552e36 ;
init_grad[ 513 ] = 36'h551c78e31 ;
init_grad[ 514 ] = 36'h54e3b2e2d ;
init_grad[ 515 ] = 36'h54aafee28 ;
init_grad[ 516 ] = 36'h54725ce23 ;
init_grad[ 517 ] = 36'h5439cee1e ;
init_grad[ 518 ] = 36'h540152e1a ;
init_grad[ 519 ] = 36'h53c8e8e15 ;
init_grad[ 520 ] = 36'h539092e10 ;
init_grad[ 521 ] = 36'h53584ee0c ;
init_grad[ 522 ] = 36'h53201ee07 ;
init_grad[ 523 ] = 36'h52e7fee02 ;
init_grad[ 524 ] = 36'h52aff2dfe ;
init_grad[ 525 ] = 36'h5277fadf9 ;
init_grad[ 526 ] = 36'h524012df5 ;
init_grad[ 527 ] = 36'h52083edf0 ;
init_grad[ 528 ] = 36'h51d07cdeb ;
init_grad[ 529 ] = 36'h5198ccde7 ;
init_grad[ 530 ] = 36'h516130de2 ;
init_grad[ 531 ] = 36'h5129a4dde ;
init_grad[ 532 ] = 36'h50f22cdd9 ;
init_grad[ 533 ] = 36'h50bac6dd5 ;
init_grad[ 534 ] = 36'h508370dd0 ;
init_grad[ 535 ] = 36'h504c2edcb ;
init_grad[ 536 ] = 36'h5014fedc7 ;
init_grad[ 537 ] = 36'h4fdde0dc2 ;
init_grad[ 538 ] = 36'h4fa6d6dbe ;
init_grad[ 539 ] = 36'h4f6fdcdb9 ;
init_grad[ 540 ] = 36'h4f38f4db5 ;
init_grad[ 541 ] = 36'h4f021edb0 ;
init_grad[ 542 ] = 36'h4ecb5adac ;
init_grad[ 543 ] = 36'h4e94a8da8 ;
init_grad[ 544 ] = 36'h4e5e08da3 ;
init_grad[ 545 ] = 36'h4e277ad9f ;
init_grad[ 546 ] = 36'h4df0fed9a ;
init_grad[ 547 ] = 36'h4dba92d96 ;
init_grad[ 548 ] = 36'h4d843ad91 ;
init_grad[ 549 ] = 36'h4d4df2d8d ;
init_grad[ 550 ] = 36'h4d17bcd89 ;
init_grad[ 551 ] = 36'h4ce198d84 ;
init_grad[ 552 ] = 36'h4cab86d80 ;
init_grad[ 553 ] = 36'h4c7586d7b ;
init_grad[ 554 ] = 36'h4c3f96d77 ;
init_grad[ 555 ] = 36'h4c09b8d73 ;
init_grad[ 556 ] = 36'h4bd3ecd6e ;
init_grad[ 557 ] = 36'h4b9e30d6a ;
init_grad[ 558 ] = 36'h4b6886d66 ;
init_grad[ 559 ] = 36'h4b32eed61 ;
init_grad[ 560 ] = 36'h4afd68d5d ;
init_grad[ 561 ] = 36'h4ac7f2d59 ;
init_grad[ 562 ] = 36'h4a928ed54 ;
init_grad[ 563 ] = 36'h4a5d3ad50 ;
init_grad[ 564 ] = 36'h4a27f8d4c ;
init_grad[ 565 ] = 36'h49f2c8d47 ;
init_grad[ 566 ] = 36'h49bda8d43 ;
init_grad[ 567 ] = 36'h49889ad3f ;
init_grad[ 568 ] = 36'h49539cd3b ;
init_grad[ 569 ] = 36'h491eb0d36 ;
init_grad[ 570 ] = 36'h48e9d4d32 ;
init_grad[ 571 ] = 36'h48b50ad2e ;
init_grad[ 572 ] = 36'h488050d2a ;
init_grad[ 573 ] = 36'h484ba8d25 ;
init_grad[ 574 ] = 36'h481710d21 ;
init_grad[ 575 ] = 36'h47e288d1d ;
init_grad[ 576 ] = 36'h47ae12d19 ;
init_grad[ 577 ] = 36'h4779acd15 ;
init_grad[ 578 ] = 36'h474558d10 ;
init_grad[ 579 ] = 36'h471114d0c ;
init_grad[ 580 ] = 36'h46dce0d08 ;
init_grad[ 581 ] = 36'h46a8bed04 ;
init_grad[ 582 ] = 36'h4674acd00 ;
init_grad[ 583 ] = 36'h4640aacfc ;
init_grad[ 584 ] = 36'h460cbacf8 ;
init_grad[ 585 ] = 36'h45d8dacf3 ;
init_grad[ 586 ] = 36'h45a50acef ;
init_grad[ 587 ] = 36'h45714aceb ;
init_grad[ 588 ] = 36'h453d9cce7 ;
init_grad[ 589 ] = 36'h4509fece3 ;
init_grad[ 590 ] = 36'h44d670cdf ;
init_grad[ 591 ] = 36'h44a2f2cdb ;
init_grad[ 592 ] = 36'h446f84cd7 ;
init_grad[ 593 ] = 36'h443c26cd3 ;
init_grad[ 594 ] = 36'h4408daccf ;
init_grad[ 595 ] = 36'h43d59eccb ;
init_grad[ 596 ] = 36'h43a270cc7 ;
init_grad[ 597 ] = 36'h436f54cc3 ;
init_grad[ 598 ] = 36'h433c48cbf ;
init_grad[ 599 ] = 36'h43094ccbb ;
init_grad[ 600 ] = 36'h42d660cb6 ;
init_grad[ 601 ] = 36'h42a384cb2 ;
init_grad[ 602 ] = 36'h4270b8cae ;
init_grad[ 603 ] = 36'h423dfccab ;
init_grad[ 604 ] = 36'h420b50ca7 ;
init_grad[ 605 ] = 36'h41d8b4ca3 ;
init_grad[ 606 ] = 36'h41a628c9f ;
init_grad[ 607 ] = 36'h4173acc9b ;
init_grad[ 608 ] = 36'h41413ec97 ;
init_grad[ 609 ] = 36'h410ee2c93 ;
init_grad[ 610 ] = 36'h40dc96c8f ;
init_grad[ 611 ] = 36'h40aa58c8b ;
init_grad[ 612 ] = 36'h40782ac87 ;
init_grad[ 613 ] = 36'h40460ec83 ;
init_grad[ 614 ] = 36'h4013fec7f ;
init_grad[ 615 ] = 36'h3fe200c7b ;
init_grad[ 616 ] = 36'h3fb012c77 ;
init_grad[ 617 ] = 36'h3f7e32c73 ;
init_grad[ 618 ] = 36'h3f4c62c70 ;
init_grad[ 619 ] = 36'h3f1aa2c6c ;
init_grad[ 620 ] = 36'h3ee8f2c68 ;
init_grad[ 621 ] = 36'h3eb750c64 ;
init_grad[ 622 ] = 36'h3e85bec60 ;
init_grad[ 623 ] = 36'h3e543cc5c ;
init_grad[ 624 ] = 36'h3e22cac58 ;
init_grad[ 625 ] = 36'h3df166c55 ;
init_grad[ 626 ] = 36'h3dc012c51 ;
init_grad[ 627 ] = 36'h3d8eccc4d ;
init_grad[ 628 ] = 36'h3d5d96c49 ;
init_grad[ 629 ] = 36'h3d2c70c45 ;
init_grad[ 630 ] = 36'h3cfb5ac42 ;
init_grad[ 631 ] = 36'h3cca50c3e ;
init_grad[ 632 ] = 36'h3c9958c3a ;
init_grad[ 633 ] = 36'h3c686ec36 ;
init_grad[ 634 ] = 36'h3c3794c32 ;
init_grad[ 635 ] = 36'h3c06c8c2f ;
init_grad[ 636 ] = 36'h3bd60cc2b ;
init_grad[ 637 ] = 36'h3ba55ec27 ;
init_grad[ 638 ] = 36'h3b74c0c23 ;
init_grad[ 639 ] = 36'h3b4430c20 ;
init_grad[ 640 ] = 36'h3b13aec1c ;
init_grad[ 641 ] = 36'h3ae33ec18 ;
init_grad[ 642 ] = 36'h3ab2dac14 ;
init_grad[ 643 ] = 36'h3a8286c11 ;
init_grad[ 644 ] = 36'h3a5242c0d ;
init_grad[ 645 ] = 36'h3a220ac09 ;
init_grad[ 646 ] = 36'h39f1e4c06 ;
init_grad[ 647 ] = 36'h39c1cac02 ;
init_grad[ 648 ] = 36'h3991c0bfe ;
init_grad[ 649 ] = 36'h3961c6bfb ;
init_grad[ 650 ] = 36'h3931d8bf7 ;
init_grad[ 651 ] = 36'h3901fabf3 ;
init_grad[ 652 ] = 36'h38d22abf0 ;
init_grad[ 653 ] = 36'h38a26abec ;
init_grad[ 654 ] = 36'h3872b8be8 ;
init_grad[ 655 ] = 36'h384314be5 ;
init_grad[ 656 ] = 36'h381380be1 ;
init_grad[ 657 ] = 36'h37e3f8bde ;
init_grad[ 658 ] = 36'h37b480bda ;
init_grad[ 659 ] = 36'h378516bd6 ;
init_grad[ 660 ] = 36'h3755babd3 ;
init_grad[ 661 ] = 36'h37266ebcf ;
init_grad[ 662 ] = 36'h36f730bcc ;
init_grad[ 663 ] = 36'h36c800bc8 ;
init_grad[ 664 ] = 36'h3698debc4 ;
init_grad[ 665 ] = 36'h3669cabc1 ;
init_grad[ 666 ] = 36'h363ac4bbd ;
init_grad[ 667 ] = 36'h360bccbba ;
init_grad[ 668 ] = 36'h35dce4bb6 ;
init_grad[ 669 ] = 36'h35ae0abb3 ;
init_grad[ 670 ] = 36'h357f3cbaf ;
init_grad[ 671 ] = 36'h35507ebac ;
init_grad[ 672 ] = 36'h3521ceba8 ;
init_grad[ 673 ] = 36'h34f32cba5 ;
init_grad[ 674 ] = 36'h34c496ba1 ;
init_grad[ 675 ] = 36'h349610b9e ;
init_grad[ 676 ] = 36'h346798b9a ;
init_grad[ 677 ] = 36'h34392eb97 ;
init_grad[ 678 ] = 36'h340ad2b93 ;
init_grad[ 679 ] = 36'h33dc84b90 ;
init_grad[ 680 ] = 36'h33ae44b8c ;
init_grad[ 681 ] = 36'h338012b89 ;
init_grad[ 682 ] = 36'h3351ecb85 ;
init_grad[ 683 ] = 36'h3323d6b82 ;
init_grad[ 684 ] = 36'h32f5ccb7e ;
init_grad[ 685 ] = 36'h32c7d2b7b ;
init_grad[ 686 ] = 36'h3299e4b77 ;
init_grad[ 687 ] = 36'h326c04b74 ;
init_grad[ 688 ] = 36'h323e32b71 ;
init_grad[ 689 ] = 36'h32106eb6d ;
init_grad[ 690 ] = 36'h31e2b8b6a ;
init_grad[ 691 ] = 36'h31b50eb66 ;
init_grad[ 692 ] = 36'h318774b63 ;
init_grad[ 693 ] = 36'h3159e6b60 ;
init_grad[ 694 ] = 36'h312c66b5c ;
init_grad[ 695 ] = 36'h30fef2b59 ;
init_grad[ 696 ] = 36'h30d18eb55 ;
init_grad[ 697 ] = 36'h30a436b52 ;
init_grad[ 698 ] = 36'h3076ecb4f ;
init_grad[ 699 ] = 36'h3049b0b4b ;
init_grad[ 700 ] = 36'h301c80b48 ;
init_grad[ 701 ] = 36'h2fef5eb45 ;
init_grad[ 702 ] = 36'h2fc24ab41 ;
init_grad[ 703 ] = 36'h2f9544b3e ;
init_grad[ 704 ] = 36'h2f684ab3b ;
init_grad[ 705 ] = 36'h2f3b5eb37 ;
init_grad[ 706 ] = 36'h2f0e7eb34 ;
init_grad[ 707 ] = 36'h2ee1acb31 ;
init_grad[ 708 ] = 36'h2eb4e8b2d ;
init_grad[ 709 ] = 36'h2e8830b2a ;
init_grad[ 710 ] = 36'h2e5b86b27 ;
init_grad[ 711 ] = 36'h2e2eeab23 ;
init_grad[ 712 ] = 36'h2e025ab20 ;
init_grad[ 713 ] = 36'h2dd5d8b1d ;
init_grad[ 714 ] = 36'h2da962b1a ;
init_grad[ 715 ] = 36'h2d7cfab16 ;
init_grad[ 716 ] = 36'h2d509eb13 ;
init_grad[ 717 ] = 36'h2d2450b10 ;
init_grad[ 718 ] = 36'h2cf80eb0d ;
init_grad[ 719 ] = 36'h2ccbdab09 ;
init_grad[ 720 ] = 36'h2c9fb2b06 ;
init_grad[ 721 ] = 36'h2c7398b03 ;
init_grad[ 722 ] = 36'h2c478ab00 ;
init_grad[ 723 ] = 36'h2c1b8aafc ;
init_grad[ 724 ] = 36'h2bef96af9 ;
init_grad[ 725 ] = 36'h2bc3b0af6 ;
init_grad[ 726 ] = 36'h2b97d6af3 ;
init_grad[ 727 ] = 36'h2b6c0aaf0 ;
init_grad[ 728 ] = 36'h2b4048aec ;
init_grad[ 729 ] = 36'h2b1496ae9 ;
init_grad[ 730 ] = 36'h2ae8eeae6 ;
init_grad[ 731 ] = 36'h2abd54ae3 ;
init_grad[ 732 ] = 36'h2a91c8ae0 ;
init_grad[ 733 ] = 36'h2a6646adc ;
init_grad[ 734 ] = 36'h2a3ad2ad9 ;
init_grad[ 735 ] = 36'h2a0f6cad6 ;
init_grad[ 736 ] = 36'h29e410ad3 ;
init_grad[ 737 ] = 36'h29b8c2ad0 ;
init_grad[ 738 ] = 36'h298d82acd ;
init_grad[ 739 ] = 36'h29624caca ;
init_grad[ 740 ] = 36'h293724ac6 ;
init_grad[ 741 ] = 36'h290c08ac3 ;
init_grad[ 742 ] = 36'h28e0f8ac0 ;
init_grad[ 743 ] = 36'h28b5f6abd ;
init_grad[ 744 ] = 36'h288b00aba ;
init_grad[ 745 ] = 36'h286016ab7 ;
init_grad[ 746 ] = 36'h283538ab4 ;
init_grad[ 747 ] = 36'h280a66ab1 ;
init_grad[ 748 ] = 36'h27dfa2aae ;
init_grad[ 749 ] = 36'h27b4eaaab ;
init_grad[ 750 ] = 36'h278a3caa7 ;
init_grad[ 751 ] = 36'h275f9eaa4 ;
init_grad[ 752 ] = 36'h27350aaa1 ;
init_grad[ 753 ] = 36'h270a82a9e ;
init_grad[ 754 ] = 36'h26e008a9b ;
init_grad[ 755 ] = 36'h26b598a98 ;
init_grad[ 756 ] = 36'h268b36a95 ;
init_grad[ 757 ] = 36'h2660e0a92 ;
init_grad[ 758 ] = 36'h263696a8f ;
init_grad[ 759 ] = 36'h260c58a8c ;
init_grad[ 760 ] = 36'h25e226a89 ;
init_grad[ 761 ] = 36'h25b800a86 ;
init_grad[ 762 ] = 36'h258de6a83 ;
init_grad[ 763 ] = 36'h2563d8a80 ;
init_grad[ 764 ] = 36'h2539d6a7d ;
init_grad[ 765 ] = 36'h250fe0a7a ;
init_grad[ 766 ] = 36'h24e5f6a77 ;
init_grad[ 767 ] = 36'h24bc18a74 ;
init_grad[ 768 ] = 36'h249248a71 ;
init_grad[ 769 ] = 36'h246882a6e ;
init_grad[ 770 ] = 36'h243ec8a6b ;
init_grad[ 771 ] = 36'h24151aa68 ;
init_grad[ 772 ] = 36'h23eb78a65 ;
init_grad[ 773 ] = 36'h23c1e2a62 ;
init_grad[ 774 ] = 36'h239856a5f ;
init_grad[ 775 ] = 36'h236ed8a5c ;
init_grad[ 776 ] = 36'h234566a59 ;
init_grad[ 777 ] = 36'h231bfea56 ;
init_grad[ 778 ] = 36'h22f2a4a53 ;
init_grad[ 779 ] = 36'h22c954a50 ;
init_grad[ 780 ] = 36'h22a010a4e ;
init_grad[ 781 ] = 36'h2276d8a4b ;
init_grad[ 782 ] = 36'h224daca48 ;
init_grad[ 783 ] = 36'h22248ca45 ;
init_grad[ 784 ] = 36'h21fb76a42 ;
init_grad[ 785 ] = 36'h21d26ca3f ;
init_grad[ 786 ] = 36'h21a96ea3c ;
init_grad[ 787 ] = 36'h21807ca39 ;
init_grad[ 788 ] = 36'h215796a36 ;
init_grad[ 789 ] = 36'h212ebaa33 ;
init_grad[ 790 ] = 36'h2105eca31 ;
init_grad[ 791 ] = 36'h20dd28a2e ;
init_grad[ 792 ] = 36'h20b46ea2b ;
init_grad[ 793 ] = 36'h208bc2a28 ;
init_grad[ 794 ] = 36'h206320a25 ;
init_grad[ 795 ] = 36'h203a8aa22 ;
init_grad[ 796 ] = 36'h201200a1f ;
init_grad[ 797 ] = 36'h1fe980a1c ;
init_grad[ 798 ] = 36'h1fc10ca1a ;
init_grad[ 799 ] = 36'h1f98a4a17 ;
init_grad[ 800 ] = 36'h1f7046a14 ;
init_grad[ 801 ] = 36'h1f47f4a11 ;
init_grad[ 802 ] = 36'h1f1faea0e ;
init_grad[ 803 ] = 36'h1ef772a0c ;
init_grad[ 804 ] = 36'h1ecf42a09 ;
init_grad[ 805 ] = 36'h1ea71ea06 ;
init_grad[ 806 ] = 36'h1e7f04a03 ;
init_grad[ 807 ] = 36'h1e56f4a00 ;
init_grad[ 808 ] = 36'h1e2ef29fe ;
init_grad[ 809 ] = 36'h1e06fa9fb ;
init_grad[ 810 ] = 36'h1ddf0c9f8 ;
init_grad[ 811 ] = 36'h1db72c9f5 ;
init_grad[ 812 ] = 36'h1d8f549f2 ;
init_grad[ 813 ] = 36'h1d678a9f0 ;
init_grad[ 814 ] = 36'h1d3fc89ed ;
init_grad[ 815 ] = 36'h1d18149ea ;
init_grad[ 816 ] = 36'h1cf0689e7 ;
init_grad[ 817 ] = 36'h1cc8ca9e5 ;
init_grad[ 818 ] = 36'h1ca1369e2 ;
init_grad[ 819 ] = 36'h1c79ac9df ;
init_grad[ 820 ] = 36'h1c522e9dc ;
init_grad[ 821 ] = 36'h1c2aba9da ;
init_grad[ 822 ] = 36'h1c03529d7 ;
init_grad[ 823 ] = 36'h1bdbf49d4 ;
init_grad[ 824 ] = 36'h1bb4a29d1 ;
init_grad[ 825 ] = 36'h1b8d5a9cf ;
init_grad[ 826 ] = 36'h1b661e9cc ;
init_grad[ 827 ] = 36'h1b3eec9c9 ;
init_grad[ 828 ] = 36'h1b17c49c7 ;
init_grad[ 829 ] = 36'h1af0a89c4 ;
init_grad[ 830 ] = 36'h1ac9969c1 ;
init_grad[ 831 ] = 36'h1aa2909be ;
init_grad[ 832 ] = 36'h1a7b949bc ;
init_grad[ 833 ] = 36'h1a54a29b9 ;
init_grad[ 834 ] = 36'h1a2dbc9b6 ;
init_grad[ 835 ] = 36'h1a06e09b4 ;
init_grad[ 836 ] = 36'h19e0109b1 ;
init_grad[ 837 ] = 36'h19b94a9ae ;
init_grad[ 838 ] = 36'h19928e9ac ;
init_grad[ 839 ] = 36'h196bdc9a9 ;
init_grad[ 840 ] = 36'h1945369a6 ;
init_grad[ 841 ] = 36'h191e9a9a4 ;
init_grad[ 842 ] = 36'h18f80a9a1 ;
init_grad[ 843 ] = 36'h18d18299f ;
init_grad[ 844 ] = 36'h18ab0699c ;
init_grad[ 845 ] = 36'h188494999 ;
init_grad[ 846 ] = 36'h185e2e997 ;
init_grad[ 847 ] = 36'h1837d2994 ;
init_grad[ 848 ] = 36'h181180991 ;
init_grad[ 849 ] = 36'h17eb3898f ;
init_grad[ 850 ] = 36'h17c4fa98c ;
init_grad[ 851 ] = 36'h179ec898a ;
init_grad[ 852 ] = 36'h1778a0987 ;
init_grad[ 853 ] = 36'h175282984 ;
init_grad[ 854 ] = 36'h172c6e982 ;
init_grad[ 855 ] = 36'h17066697f ;
init_grad[ 856 ] = 36'h16e06697d ;
init_grad[ 857 ] = 36'h16ba7297a ;
init_grad[ 858 ] = 36'h169488977 ;
init_grad[ 859 ] = 36'h166ea8975 ;
init_grad[ 860 ] = 36'h1648d4972 ;
init_grad[ 861 ] = 36'h162308970 ;
init_grad[ 862 ] = 36'h15fd4896d ;
init_grad[ 863 ] = 36'h15d79096b ;
init_grad[ 864 ] = 36'h15b1e4968 ;
init_grad[ 865 ] = 36'h158c42966 ;
init_grad[ 866 ] = 36'h1566aa963 ;
init_grad[ 867 ] = 36'h15411c960 ;
init_grad[ 868 ] = 36'h151b9895e ;
init_grad[ 869 ] = 36'h14f61e95b ;
init_grad[ 870 ] = 36'h14d0b0959 ;
init_grad[ 871 ] = 36'h14ab4a956 ;
init_grad[ 872 ] = 36'h1485f0954 ;
init_grad[ 873 ] = 36'h14609e951 ;
init_grad[ 874 ] = 36'h143b5694f ;
init_grad[ 875 ] = 36'h14161a94c ;
init_grad[ 876 ] = 36'h13f0e694a ;
init_grad[ 877 ] = 36'h13cbbe947 ;
init_grad[ 878 ] = 36'h13a6a0945 ;
init_grad[ 879 ] = 36'h13818a942 ;
init_grad[ 880 ] = 36'h135c80940 ;
init_grad[ 881 ] = 36'h13377e93d ;
init_grad[ 882 ] = 36'h13128893b ;
init_grad[ 883 ] = 36'h12ed9a938 ;
init_grad[ 884 ] = 36'h12c8b6936 ;
init_grad[ 885 ] = 36'h12a3de933 ;
init_grad[ 886 ] = 36'h127f0e931 ;
init_grad[ 887 ] = 36'h125a4892e ;
init_grad[ 888 ] = 36'h12358c92c ;
init_grad[ 889 ] = 36'h1210da92a ;
init_grad[ 890 ] = 36'h11ec32927 ;
init_grad[ 891 ] = 36'h11c794925 ;
init_grad[ 892 ] = 36'h11a300922 ;
init_grad[ 893 ] = 36'h117e76920 ;
init_grad[ 894 ] = 36'h1159f491d ;
init_grad[ 895 ] = 36'h11357c91b ;
init_grad[ 896 ] = 36'h111110918 ;
init_grad[ 897 ] = 36'h10ecac916 ;
init_grad[ 898 ] = 36'h10c852914 ;
init_grad[ 899 ] = 36'h10a400911 ;
init_grad[ 900 ] = 36'h107fba90f ;
init_grad[ 901 ] = 36'h105b7c90c ;
init_grad[ 902 ] = 36'h10374a90a ;
init_grad[ 903 ] = 36'h101320908 ;
init_grad[ 904 ] = 36'hfef00905 ;
init_grad[ 905 ] = 36'hfcae8903 ;
init_grad[ 906 ] = 36'hfa6dc900 ;
init_grad[ 907 ] = 36'hf82d88fe ;
init_grad[ 908 ] = 36'hf5ede8fc ;
init_grad[ 909 ] = 36'hf3aee8f9 ;
init_grad[ 910 ] = 36'hf17068f7 ;
init_grad[ 911 ] = 36'hef3288f4 ;
init_grad[ 912 ] = 36'hecf548f2 ;
init_grad[ 913 ] = 36'heab8a8f0 ;
init_grad[ 914 ] = 36'he87ca8ed ;
init_grad[ 915 ] = 36'he64128eb ;
init_grad[ 916 ] = 36'he40648e9 ;
init_grad[ 917 ] = 36'he1cbe8e6 ;
init_grad[ 918 ] = 36'hdf9248e4 ;
init_grad[ 919 ] = 36'hdd5928e2 ;
init_grad[ 920 ] = 36'hdb2088df ;
init_grad[ 921 ] = 36'hd8e8a8dd ;
init_grad[ 922 ] = 36'hd6b148db ;
init_grad[ 923 ] = 36'hd47a68d8 ;
init_grad[ 924 ] = 36'hd24448d6 ;
init_grad[ 925 ] = 36'hd00ea8d4 ;
init_grad[ 926 ] = 36'hcdd988d1 ;
init_grad[ 927 ] = 36'hcba528cf ;
init_grad[ 928 ] = 36'hc97148cd ;
init_grad[ 929 ] = 36'hc73de8ca ;
init_grad[ 930 ] = 36'hc50b28c8 ;
init_grad[ 931 ] = 36'hc2d908c6 ;
init_grad[ 932 ] = 36'hc0a768c4 ;
init_grad[ 933 ] = 36'hbe7668c1 ;
init_grad[ 934 ] = 36'hbc4608bf ;
init_grad[ 935 ] = 36'hba1628bd ;
init_grad[ 936 ] = 36'hb7e6c8ba ;
init_grad[ 937 ] = 36'hb5b828b8 ;
init_grad[ 938 ] = 36'hb389e8b6 ;
init_grad[ 939 ] = 36'hb15c68b4 ;
init_grad[ 940 ] = 36'haf2f68b1 ;
init_grad[ 941 ] = 36'had02e8af ;
init_grad[ 942 ] = 36'haad708ad ;
init_grad[ 943 ] = 36'ha8aba8ab ;
init_grad[ 944 ] = 36'ha680e8a8 ;
init_grad[ 945 ] = 36'ha456c8a6 ;
init_grad[ 946 ] = 36'ha22d28a4 ;
init_grad[ 947 ] = 36'ha00408a2 ;
init_grad[ 948 ] = 36'h9ddb889f ;
init_grad[ 949 ] = 36'h9bb3a89d ;
init_grad[ 950 ] = 36'h998c489b ;
init_grad[ 951 ] = 36'h97656899 ;
init_grad[ 952 ] = 36'h953f2896 ;
init_grad[ 953 ] = 36'h93196894 ;
init_grad[ 954 ] = 36'h90f44892 ;
init_grad[ 955 ] = 36'h8ecfa890 ;
init_grad[ 956 ] = 36'h8caba88d ;
init_grad[ 957 ] = 36'h8a88288b ;
init_grad[ 958 ] = 36'h88652889 ;
init_grad[ 959 ] = 36'h8642c887 ;
init_grad[ 960 ] = 36'h8420e885 ;
init_grad[ 961 ] = 36'h81ffa882 ;
init_grad[ 962 ] = 36'h7fdee880 ;
init_grad[ 963 ] = 36'h7dbec87e ;
init_grad[ 964 ] = 36'h7b9f087c ;
init_grad[ 965 ] = 36'h7980087a ;
init_grad[ 966 ] = 36'h77616878 ;
init_grad[ 967 ] = 36'h75436875 ;
init_grad[ 968 ] = 36'h7325e873 ;
init_grad[ 969 ] = 36'h71090871 ;
init_grad[ 970 ] = 36'h6eeca86f ;
init_grad[ 971 ] = 36'h6cd0c86d ;
init_grad[ 972 ] = 36'h6ab5886b ;
init_grad[ 973 ] = 36'h689ac868 ;
init_grad[ 974 ] = 36'h66808866 ;
init_grad[ 975 ] = 36'h6466e864 ;
init_grad[ 976 ] = 36'h624dc862 ;
init_grad[ 977 ] = 36'h60352860 ;
init_grad[ 978 ] = 36'h5e1d085e ;
init_grad[ 979 ] = 36'h5c05885b ;
init_grad[ 980 ] = 36'h59ee8859 ;
init_grad[ 981 ] = 36'h57d80857 ;
init_grad[ 982 ] = 36'h55c22855 ;
init_grad[ 983 ] = 36'h53acc853 ;
init_grad[ 984 ] = 36'h5197e851 ;
init_grad[ 985 ] = 36'h4f83884f ;
init_grad[ 986 ] = 36'h4d6fc84d ;
init_grad[ 987 ] = 36'h4b5c884b ;
init_grad[ 988 ] = 36'h4949c848 ;
init_grad[ 989 ] = 36'h47378846 ;
init_grad[ 990 ] = 36'h4525c844 ;
init_grad[ 991 ] = 36'h4314a842 ;
init_grad[ 992 ] = 36'h41040840 ;
init_grad[ 993 ] = 36'h3ef3e83e ;
init_grad[ 994 ] = 36'h3ce4483c ;
init_grad[ 995 ] = 36'h3ad5283a ;
init_grad[ 996 ] = 36'h38c6a838 ;
init_grad[ 997 ] = 36'h36b8a836 ;
init_grad[ 998 ] = 36'h34ab2833 ;
init_grad[ 999 ] = 36'h329e2831 ;
init_grad[ 1000 ] = 36'h3091a82f ;
init_grad[ 1001 ] = 36'h2e85a82d ;
init_grad[ 1002 ] = 36'h2c7a482b ;
init_grad[ 1003 ] = 36'h2a6f4829 ;
init_grad[ 1004 ] = 36'h2864e827 ;
init_grad[ 1005 ] = 36'h265b0825 ;
init_grad[ 1006 ] = 36'h2451a823 ;
init_grad[ 1007 ] = 36'h2248c821 ;
init_grad[ 1008 ] = 36'h2040681f ;
init_grad[ 1009 ] = 36'h1e38881d ;
init_grad[ 1010 ] = 36'h1c31481b ;
init_grad[ 1011 ] = 36'h1a2a6819 ;
init_grad[ 1012 ] = 36'h18242817 ;
init_grad[ 1013 ] = 36'h161e4815 ;
init_grad[ 1014 ] = 36'h14190813 ;
init_grad[ 1015 ] = 36'h12144811 ;
init_grad[ 1016 ] = 36'h1010080f ;
init_grad[ 1017 ] = 36'he0c480d ;
init_grad[ 1018 ] = 36'hc08e80b ;
init_grad[ 1019 ] = 36'ha062809 ;
init_grad[ 1020 ] = 36'h803e807 ;
init_grad[ 1021 ] = 36'h6022804 ;
init_grad[ 1022 ] = 36'h400e802 ;
init_grad[ 1023 ] = 36'h2002800 ;

    end


endmodule