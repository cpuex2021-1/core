module tx(
    input wire clk,rst,
    input wire [7:0] dout,
    input wire 
);

endmodule