`timescale 1ns / 1ps
import axi_vip_pkg::*;
import design_2_axi_vip_0_0_pkg::*;


module simtop();
    logic clk, rst;
    logic rxd, txd;
    logic [15:0] LED;
    parameter STEP = 50; // clk(#10) * 5
    logic [31:0] count;

    task uart(input logic [7:0] data);
    begin
    #STEP rxd = 0;
    #STEP rxd = data[0];
    #STEP rxd = data[1];
    #STEP rxd = data[2];
    #STEP rxd = data[3];
    #STEP rxd = data[4];
    #STEP rxd = data[5];
    #STEP rxd = data[6];
    #STEP rxd = data[7];
    #STEP rxd = 1;
    end
    endtask
    always  begin
        clk = 1'b0;
        #5 clk = 1'b1;
        #5 count = count+1;
    end

        logic [7:0] data;
/*logic [7:0] contest_bin [0:1299] = {
  8'h00, 8'h00, 8'h8c, 8'hc2, 8'h00, 8'h00, 8'h0c, 8'h42, 8'h00, 8'h00, 8'ha0, 8'hc1,
  8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'hf0, 8'h41, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h48, 8'h42, 8'h00, 8'h00, 8'h48, 8'h42, 8'h00, 8'h00, 8'h7f, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'ha0, 8'h41,
  8'h00, 8'h00, 8'h82, 8'h42, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h41,
  8'h00, 8'h00, 8'h34, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h52, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc8, 8'h41,
  8'h00, 8'h00, 8'h20, 8'h42, 8'h00, 8'h00, 8'h8c, 8'h42, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43,
  8'h00, 8'h00, 8'h52, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hf0, 8'h41, 8'h00, 8'h00, 8'hf0, 8'h41,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h80, 8'hbf, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'h20, 8'h41,
  8'h00, 8'h00, 8'hf0, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hc1,
  8'h00, 8'h00, 8'ha0, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'hc0, 8'hbf, 8'h00, 8'h00, 8'h80, 8'hbf, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43,
  8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'hb0, 8'h41, 8'h00, 8'h00, 8'he0, 8'h41, 8'h00, 8'h00, 8'he0, 8'h41,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h42, 8'h00, 8'h00, 8'he0, 8'h41,
  8'h00, 8'h00, 8'he0, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'hc0,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h43,
  8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h70, 8'h41, 8'h00, 8'h00, 8'h70, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'ha0, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'hbf,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h70, 8'h41, 8'h00, 8'h00, 8'hc8, 8'h41, 8'h00, 8'h00, 8'hc8, 8'h41,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'hc0, 8'h00, 8'h00, 8'h8c, 8'h42,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43,
  8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h40, 8'h00, 8'h00, 8'h30, 8'h41,
  8'h00, 8'h00, 8'h34, 8'h42, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'h42,
  8'h00, 8'h00, 8'h20, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hf0, 8'h41,
  8'h00, 8'h00, 8'h34, 8'h42, 8'h00, 8'h00, 8'h96, 8'h42, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'hc8, 8'h41, 8'h00, 8'h00, 8'h24, 8'h42, 8'h00, 8'h00, 8'h8c, 8'h42,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h40, 8'h00, 8'h00, 8'h20, 8'h42,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc8, 8'h42, 8'h00, 8'h00, 8'ha0, 8'h40,
  8'h00, 8'h00, 8'h48, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0c, 8'hc2,
  8'h00, 8'h00, 8'h16, 8'h43, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h48, 8'h43, 8'h00, 8'h00, 8'h48, 8'h43,
  8'h00, 8'h00, 8'h48, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hc8, 8'h41,
  8'h00, 8'h00, 8'h20, 8'h41, 8'h00, 8'h00, 8'h20, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'ha0, 8'hc0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h7a, 8'h43, 8'h00, 8'h00, 8'h53, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h00, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h03, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'hc8, 8'h41, 8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'ha0, 8'h41,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h8c, 8'h42,
  8'h00, 8'h00, 8'h80, 8'h3f, 8'h9a, 8'h99, 8'h99, 8'h3e, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7f, 8'h43,
  8'h02, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'ha0, 8'h41,
  8'h00, 8'h00, 8'ha0, 8'h41, 8'h00, 8'h00, 8'hc8, 8'h42, 8'h00, 8'h00, 8'h20, 8'h42,
  8'h00, 8'h00, 8'hf0, 8'h42, 8'h00, 8'h00, 8'h80, 8'h3f, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'h00, 8'h00, 8'h16, 8'h43, 8'h00, 8'h00, 8'h7f, 8'h43, 8'h00, 8'h00, 8'h7f, 8'h43,
  8'h00, 8'h00, 8'h7f, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00,
  8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'hbf, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h43, 8'h00, 8'h00, 8'h80, 8'h3f,
  8'hcd, 8'hcc, 8'h4c, 8'h3e, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7f, 8'h43,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00,
  8'hff, 8'hff, 8'hff, 8'hff, 8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00,
  8'h04, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h05, 8'h00, 8'h00, 8'h00,
  8'h06, 8'h00, 8'h00, 8'h00, 8'h07, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'h08, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h09, 8'h00, 8'h00, 8'h00,
  8'h0a, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h0c, 8'h00, 8'h00, 8'h00,
  8'hff, 8'hff, 8'hff, 8'hff, 8'h0d, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'h0e, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff, 8'h0f, 8'h00, 8'h00, 8'h00,
  8'hff, 8'hff, 8'hff, 8'hff, 8'h10, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'hff, 8'hff, 8'hff, 8'hff, 8'h0b, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
  8'h01, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00,
  8'h04, 8'h00, 8'h00, 8'h00, 8'h06, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'h63, 8'h00, 8'h00, 8'h00, 8'h09, 8'h00, 8'h00, 8'h00, 8'h08, 8'h00, 8'h00, 8'h00,
  8'h07, 8'h00, 8'h00, 8'h00, 8'h05, 8'h00, 8'h00, 8'h00, 8'hff, 8'hff, 8'hff, 8'hff,
  8'hff, 8'hff, 8'hff, 8'hff
};*/
logic [7:0] send_bin[0:167] = {
  8'h15, 8'h00, 8'h40, 8'h00, 8'h84, 8'h0a, 8'h40, 8'h08, 8'h04, 8'h0c, 8'hc0, 8'h01,
  8'h04, 8'h08, 8'h00, 8'h02, 8'h84, 8'h02, 8'h40, 8'h02, 8'h04, 8'h14, 8'h80, 8'h01,
  8'hb6, 8'h01, 8'h00, 8'h00, 8'hc4, 8'h0c, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00,
  8'h76, 8'h02, 8'h00, 8'h00, 8'h44, 8'h0c, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00,
  8'h84, 8'h0c, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00, 8'h04, 8'h0e, 8'h80, 8'h01,
  8'hb6, 8'h01, 8'h00, 8'h00, 8'h36, 8'h02, 8'h00, 8'h00, 8'h44, 8'h0c, 8'h80, 8'h01,
  8'hb6, 8'h01, 8'h00, 8'h00, 8'h84, 8'h0c, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00,
  8'h04, 8'h0e, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00, 8'h36, 8'h02, 8'h00, 8'h00,
  8'h84, 8'h0c, 8'h80, 8'h01, 8'hb6, 8'h01, 8'h00, 8'h00, 8'h44, 8'h0d, 8'h80, 8'h01,
  8'hb6, 8'h01, 8'h00, 8'h00, 8'hb6, 8'h01, 8'h00, 8'h00, 8'h76, 8'h02, 8'h00, 8'h00,
  8'h04, 8'h00, 8'h90, 8'h01, 8'h04, 8'h0c, 8'hc0, 8'h01, 8'h04, 8'h08, 8'h00, 8'h02,
  8'h84, 8'h02, 8'h40, 8'h02, 8'hf6, 8'h01, 8'h00, 8'h00, 8'h36, 8'h02, 8'h00, 8'h00,
  8'hf6, 8'h01, 8'h00, 8'h00, 8'h36, 8'h02, 8'h00, 8'h00, 8'hf6, 8'h01, 8'h00, 8'h00,
  8'h76, 8'h02, 8'h00, 8'h00, 8'hc4, 8'hff, 8'hbf, 8'h31, 8'h0e, 8'hc8, 8'hff, 8'h37
};

        int i;
    initial begin
        rxd = 1;
        rst = 1'b0;
        
        #13 rst = 1'b1;  
        count = -33;      
        //repeat(30) 
        #500;
        //uart(12);
        //uart(0);
        //uart(0);
        //uart(0);
        
        //uart(8'd5);
        //uart(0);
        //uart(8'd128);
        //uart(1);
        
        //uart(182);
        //uart(1);
        //uart(0);
        //uart(0);
        
        //uart(135);
        //uart(0);
        //uart(0);
        //uart(0);
        
        //uart(0);
        /*for(i=0; i<1300; i=i+1) begin
            uart(contest_bin[i]);
        end*/
        uart(168);
        uart(0);
        uart(0);
        uart(0);
        
        
        for(i=0; i<168; i=i+1) begin
            uart(send_bin[i]);
        end
        //end
                
    end

    design_2_wrapper dut(.sys_clock (clk), .reset (rst), .rxd(rxd), .txd(txd), .LED);
    design_2_axi_vip_0_0_slv_mem_t agent;
    initial begin

       agent = new("AXI Slave Agent", dut.design_2_i.axi_vip_0.inst.IF);
        agent.start_slave();
    end
endmodule