typedef struct {
    logic AXI_RADDR;
} axi;